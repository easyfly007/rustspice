* RC Lowpass Filter for AC Analysis Test
* Cutoff frequency fc = 1/(2*pi*R*C) = 1/(2*pi*1k*1u) = 159.15 Hz

V1 in 0 DC 0 AC 1 0
R1 in out 1k
C1 out 0 1u

.ac dec 10 1 1meg
.end
